`timescale 1ns / 1ps

module wbuffer_tb();

endmodule