`timescale 1ns / 1ps

module wbuffer_tb();

    wire [4:0] a[2:0];
endmodule